library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.all;

entity MUL_DIV_MOD is
	port (
	);
end MUL_DIV_MOD;

architecture Behavioural of MUL_DIV_MOD is
begin
end Behavioural;


